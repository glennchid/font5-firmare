`define SIM_MODE

