//`define INCLUDE_TESTBENCH

//`define DOUBLE_CONTROL_REGS

//`define ADDPIPEREGS

`define DISABLE_AUXOUTS

//`define LOAD_ATF_DEFAULTS